LIBRARY IEEE; -- These lines informs the compiler that the library IEEE is used
USE IEEE.std_logic_1164.all; -- contains the definition for the std_logic type plus some useful conversion functions

ENTITY tb_data_bus IS END tb_data_bus;

ARCHITECTURE test of tb_data_bus IS
COMPONENT data_bus IS
PORT(data_in: IN STD_LOGIC_VECTOR(3 DOWNTO 0);        --data bus
    data_out: OUT STD_LOGIC_VECTOR(3 DOWNTO 0):="ZZZZ";
    rd_wr, clk, rst, addr: IN STD_LOGIC);                     --register read-write select, clock, register select
END COMPONENT;

SIGNAL data_in, data_out: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL clk, rst: STD_LOGIC:='0';
SIGNAL rd_wr, addr: STD_LOGIC;

BEGIN
T1: data_bus PORT MAP(data_in, data_out, rd_wr, clk, rst, addr);

data_in<="0011",
          "1010" AFTER 10 ns;

rd_wr<='1',
       '0' AFTER 20 ns;

addr<='0',
      '1' AFTER 10 ns,
      '0' AFTER 20 ns,
      '1' AFTER 30 ns;

rst<='1' AFTER 25 ns;
clk<=NOT(clk) AFTER 5 ns;
END test;
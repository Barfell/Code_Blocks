LIBRARY IEEE; -- These lines informs the compiler that the library IEEE is used
USE IEEE.std_logic_1164.all; -- contains the definition for the std_logic type plus some useful conversion functions

ENTITY tb_mux_2x1 IS END tb_mux_2x1;

ARCHITECTURE test OF tb_mux_2x1 IS
COMPONENT mux_2x1 IS
    PORT(a, b, ctrl: IN STD_LOGIC;
	q: OUT STD_LOGIC);
END COMPONENT;

SIGNAL i1: STD_LOGIC:='0';
SIGNAL i2: STD_LOGIC:='1';
SIGNAL address, result: STD_LOGIC;
BEGIN
     T1: mux_2x1 PORT MAP(a=>i1, b=>i2, ctrl=>address, q=>result);
	address<='0',
	         '1' AFTER 20 ns;
	i1<='1' AFTER 30 ns;
	i2<='0' AFTER 30 ns;
END test;